`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

module maincore(
    input clk,	//100MHz clk in
    input rst_n, //active low reset
    output[7:0] led, //status LEDss
    input usb_rx, //USB RX
    output usb_tx, //USB TX
	output led_en, led_pwm, //LED enable and PWM control for screen backlight
	//lvds outputs
	output clkout_p, clkout_n,
	output [2:0] dataout_p, dataout_n  // lvds channel 1 data outputs
	);

parameter screnn_width = 1366; //1366
parameter screnn_height = 768;  //768

parameter frame_width = 1540; //1540
parameter frame_height = 780; //780

parameter BlankingVertical = 12;
parameter BlankingHorizontal = 174;

// Total horizontal blank time is 174 pixels
parameter FrontPorchHorizontal = 30;
parameter BackPorchHorizontal = 30;
parameter hsync_pulse_size = 114;

// Total vertical blank time is 12 lines
parameter FrontPorchVertical = 3;
parameter BackPorchVertical = 4;
parameter vsync_pulse_size = 5;

parameter sync_on = 1;
parameter sync_off = ~sync_on; 

parameter integer     D = 3 ;				// Set the number of outputs per channel to be 3
parameter integer     N = 1 ;				// Set the number of channels to be 1

wire clk100_g;
wire clk72_g;
wire pixel_clk;

wire rst;

assign rst = ~rst_n;
	
assign led = rst ? 8'hAA : 8'h55; // debugging pattern
assign usb_tx = usb_rx;

reg [5:0] Red = 0;
reg [5:0] Blue = 0;
reg [5:0] Green = 0;

wire [20:0] VideoData;
wire txclk ;			
wire txclk_div ;			
wire not_tx_mmcm_lckd ;	
wire tx_mmcm_lckd ;

reg hsync = sync_off;
reg vsync = sync_off;
reg DataEnable = 0;


reg [10:0] pos_x = 0;
reg [10:0] pos_y = 0;

assign led_en = 1;
assign led_pwm = 1;

// Input Clock Buffer
BUFG bg_ref (
    .I		(clk),
    .O      (clk100_g)
	);

// Pixel Clock Generator
clk_wiz_pixel clk_pixel(
    .clk_in(clk100_g),
    .clk_out(clk72_g),
    .reset(rst)
	);

assign VideoData[20:18] = {hsync, vsync, DataEnable}; // Move to higher bits
assign VideoData[17:0]  = {Green[5:0], Red[5:0], Blue[5:0]};

// Clock Input

clock_generator_pll_7_to_1_diff_ddr #(
	.PIXEL_CLOCK		("BUF_G"),
	.INTER_CLOCK 		("BUF_G"),
	.TX_CLOCK			("BUF_G"),
	.USE_PLL			("FALSE"),
	.MMCM_MODE			(2),				// Parameter to set multiplier for MMCM to get VCO in correct operating range. 1 multiplies input clock by 7, 2 multiplies clock by 14, etc
	.CLKIN_PERIOD 		(13.889))
clkgen (                        
	.reset			(rst),
	.clkin		    (clk72_g),
	.txclk			(txclk),
	.txclk_div		(txclk_div),
	.pixel_clk		(pixel_clk),
	.status			(),
	.mmcm_lckd		(tx_mmcm_lckd)) ;

assign not_tx_mmcm_lckd = ~tx_mmcm_lckd ;

// Transmitter Logic for N D-bit channels
n_x_serdes_7_to_1_diff_ddr #(
      	.D			(D),
      	.N			(N),				// 1 channel
	.DATA_FORMAT 	("PER_CLOCK")) 			// PER_CLOCK or PER_CHANL data formatting
dataout (                      
	.dataout_p  	(dataout_p),
	.dataout_n  	(dataout_n),
	.clkout_p  		(clkout_p),
	.clkout_n  		(clkout_n),
	.txclk    		(txclk),
	.txclk_div    	(txclk_div),
	.pixel_clk		(pixel_clk),
	.reset   		(not_tx_mmcm_lckd),
	.clk_pattern  	(7'b1100011),			// Transmit a constant to make the clock
	.datain  		(VideoData)
	);



//Cycle Generator
always @(posedge pixel_clk)
begin
			// Increment horizontal position
			pos_x <= pos_x + 1;
			
			// Start horizontal blanking
			if (pos_x == screnn_width) begin
				DataEnable <= 0;
			end
			
			// Start horizontal sync
			if (pos_x == screnn_width + FrontPorchHorizontal) begin
				hsync <= sync_on;
			end
			// End horizontal sync
			else if (pos_x == screnn_width + FrontPorchHorizontal + hsync_pulse_size) begin
				hsync <= sync_off;
			end
					
			// End of line						
			if(pos_x == frame_width) begin
			        pos_x <= 0;
					pos_y <= pos_y + 1'b1;

        			// Start vertical blanking
					if(pos_y == screnn_height) begin
							DataEnable	<= 0;
					end
					
					// Start vertical sync
					if(pos_y == screnn_height + FrontPorchVertical)	begin
							vsync <= sync_on;
					end

					// End vertical sync
					if(pos_y == screnn_height + FrontPorchVertical + vsync_pulse_size) begin
							vsync <= sync_off;
					end

					// End of frame
					if(pos_y == (screnn_height + BlankingVertical)) begin
							pos_y <= 0;
							vsync <= sync_off;
					end
           end
		   else if (pos_x == 0 && pos_y < screnn_height) begin
				DataEnable <= 1;
		   end             
end

//Video Generator
always @(posedge pixel_clk)
begin
    if (DataEnable) begin
		if (pos_y < screnn_height / 2) begin
			// Generate stripes based on the horizontal position (pos_x)
			if (pos_x < screnn_width / 4) begin
				// Red stripe
				Red   <= 63;  // Maximum red
				Green <= 0;   // No green
				Blue  <= 0;   // No blue
			end else if (pos_x < screnn_width / 2) begin
				// Green stripe
				Red   <= 0;   // No red
				Green <= 63;  // Maximum green
				Blue  <= 0;   // No blue
			end else if (pos_x < 3 * screnn_width / 4) begin
				// Blue stripe
				Red   <= 0;   // No red
				Green <= 0;   // No green
				Blue  <= 63;  // Maximum blue
			end else begin
				// White stripe
				Red   <= 0;  // Maximum red
				Green <= 0;  // Maximum green
				Blue  <= 0;  // Maximum blue
			end
		end else begin
			Red   <= 0;  // No red
			Green <= 0;  // No green
			Blue  <= 0;  // No blue
		end
    end else begin
        // Blank when data enable is off
        Red   <= 0;
        Green <= 0;
        Blue  <= 0;
    end
end

endmodule